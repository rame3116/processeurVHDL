--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:03:00 05/29/2019
-- Design Name:   
-- Module Name:   /home/rahmoun/Projet_systeme_info/TestProcesseur.vhd
-- Project Name:  Projet_systeme_info
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Processeur
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TestProcesseur IS
END TestProcesseur;
 
ARCHITECTURE behavior OF TestProcesseur IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Processeur
    PORT(
         Instruction : IN  std_logic_vector(31 downto 0);
         RESET : IN  std_logic;
         CLOCK : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal Instruction : std_logic_vector(31 downto 0) := (others => '0');
   signal RESET : std_logic := '1';
   signal CLOCK : std_logic := '0';

   -- Clock period definitions
   constant CLOCK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Processeur PORT MAP (
          Instruction => Instruction,
          RESET => RESET,
          CLOCK => CLOCK
        );

   -- Clock process definitions
   CLOCK_process :process
   begin
		CLOCK <= '0';
		wait for CLOCK_period/2;
		CLOCK <= '1';
		wait for CLOCK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for CLOCK_period*10;

      -- insert stimulus here 
		Instruction <= x"61000400"; -- 6=> AFC
      wait for CLOCK_period*10;
		
		Instruction <= x"62000700";
      wait for CLOCK_period*10;
		
		Instruction <= x"55200000"; --5=> Copie
      wait for CLOCK_period*10;
		
		Instruction <= x"13120000"; --1 => Add
		wait for CLOCK_period*10;
		
--		Instruction <= x"33210000";--3=> soustraction
	--	wait for CLOCK_period*10;
		
		--Instruction <= x"24310000";--2=> multiplication
		--wait for CLOCK_period*10;
		
		Instruction <= x"80c20000"; --8 => Store à l'adresse 0c la valeur du registre 2
		wait for CLOCK_period*10;
		
		Instruction <= x"790c0000"; --7 => Load R9 @oc
		wait for CLOCK_period*10;
      wait;
   end process;

END;
